`ifndef I2C_TRANS_SVH
`define I2C_TRANS_SVH
class I2cTrans;
	byte cmd;
	byte addr;
	byte data;
endclass
`endif
