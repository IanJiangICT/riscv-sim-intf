`include "iu_seq_hello.sv"
`include "iu_seq_sim.sv"
