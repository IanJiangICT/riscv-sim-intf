`include "iu_seq_hello.sv"
