package sc_cfg;

	parameter DEC_INSN_STREAM_CAP = 272;
	parameter DEC_INSN_LIST_CAP = 16;

endpackage
